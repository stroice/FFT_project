--Delay.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;


entity Delay is
	generic(	
	  WL: integer:= 8;			-- Word Length
	  BL: integer:= 64);		   -- Buffer Length
	port(
	  rst:  in  std_logic;
	  clk:  in  std_logic;
	  Din:  in  std_logic_vector(WL -1 downto 0); 
	  Dout: out std_logic_vector(WL -1 downto 0));
end Delay;

architecture arch of Delay is

   -- At and under this limit, the delay is generated using registers. 
   -- Over this limit, the delay is generated using memories.
   constant LimitReg: integer:= 2;  

   component DelayReg 
      generic(	
         WL: integer:=8;		
         BL: integer:= 1024);		
      port(
         clk:  in  std_logic;
         Din:  in  std_logic_vector(WL -1 downto 0); 
         Dout: out std_logic_vector(WL -1 downto 0));
   end component;
   
   component DelayMem
      generic(   
        WL: integer:= 8;        
        BL: integer:= 4);        
      port(
        rst:  in  std_logic;
        clk:  in  std_logic;
        Din:  in  std_logic_vector(WL -1 downto 0); 
        Dout: out std_logic_vector(WL -1 downto 0));
   end component;

begin 

   NoDelay: if BL = 0 generate   
         Dout <= Din;
   end generate;
   
   -- At and under LimitReg, the delay is generated by using registers.
   GenReg: if (BL <= LimitReg) AND (BL > 0) generate
   
      RegBuffer: DelayReg
         generic map(	
            WL => WL,   
            BL => BL)		            
         port map(
            clk  => clk,
            Din  => Din, 
            Dout => Dout);
   
   end generate;
   
   -- Over LimitReg, the delay is generated using memories.
   GenMem: if BL > LimitReg generate
   
      MemBuffer: DelayMem
         generic map(   
            WL => WL,   
            BL => BL)                  
         port map(
            rst  => rst,
            clk  => clk,
            Din  => Din, 
            Dout => Dout);
      
   end generate;
      
end arch;
